`timescale 1 ns/1 ns


module tb_codelen_tree_build();

//localparam BITSTREAMLEN = 104;  // a fixed huffman stream
//logic [BITSTREAMLEN-1:0] bitstream = 'b11000110000111111111001100000011000000000100001011111111100110000000000011001000011011111100000010111111;

localparam BITSTREAMLEN = 100071;  // a dynamic huffman stream
logic [BITSTREAMLEN-1:0] bitstream = 'b001101111011111111101110000110010010010011101111101011100111101111010001111111100111110110101000010111010101110011100001100100111001111001100110111011100110110011100111001000011010000000001101000100111000100100100000110000000100000011001100101000101000110000011001010100010110110110100100110010101111000110100110100010100101110101011111100100111110101101001101101001101101101011101111010111111110111010110100111001101100101100101010000001010001100110000011001110011001001010000001001000001001001000001000100111101100111001110001110011011101110010011100111001010111001110011101010000111110111101111111100010101010101110111100101111001101000000000001010010111010110100100110110100011000010111110011110011110011000001100110000011001100110010111011110010111101101110101010101011110110101110011100111101111001111011110011110111100010000100101001010010100100101100110001011001100010110011000101100110001111110010100000100001010010110011111011010000010110011000101100110001011001100010110010000000110101011001100010110011000101100110001011001100010110010000000110101011001100010110011000101100110001011001000000011010101100110001011001100010110011000101100110001011001000000011010101100110001011001100011111100111111101000011011011100011100001110101011101000111101000100111100110011101100011111011000001001010101001011010100101100111110110000100111111101110001010000101101011001111101101000001011001100010110011000111111101110111110001111001101111010110111001001001111100100111110100111111001001001001000101101001101000000110101011010001110100100011110110100110111011111111110000000010100010000101011111010100100000011011001101101101100101000110100011010001000111000111000111000000000000010000100001000000101100101100101100001111110111111011111100010100010100110101101001111100100010100101010010101001000101010110101011010101000110000110000110000001111110111111011111110101111111101111101110001110001110000101001010100101010010000110110110110110111111010100011110001110101100011111000110001010101010101010100101001010100101010010000101000101000101000010000011000001100000111010111011110011101101100101100101100100101001010100101010010001110110011010000011000000010000100001000001000000100000010000000001000010000100000010101010101010101000100001000010001010111111111001100100101001010010010101011010101101010100011100011100011100000101110101110101110001001010010100111110101010111110011100000000000010101010101010110001000001100000110000000010101011010101101010100010111010111010111000101010101010101011011001000000011010101100110001011001100011111100100101001000100110010100101001110001111111001011111110001011111010000001111010000111010111111001111001111000111111011011011011011000111001011110011001111001111001101111101011110011100010000110110010101101101101110001111010100011111101110111001110110011101100111000111111111000111111111100011111111110010001001101100110110011100000000100100000001000001000100100010010000110011011100111011100111011100100111100001011110000101111000001001100000011000000110000000001101001101001101000111100100111110010011111100111000111101000011110100001111010000001111000100111100010011110001000011110110111111101101111111011011000000000001100010111000101110001100011110010111111001011111100101100111010101111010101111010101001010000101000010100010010001001000100100001100110111100110111100110111100001111000000111100000011110000000010111010101110101011100100111110011101111100111011111001111001111001111111100111111110011110011110001001111000100111100010000110000111100001111011000100111111101000111111101000111110001100010010001001000100100000111111011011111111011011111111110010100100100010010001001000101011111110101100001111010010111101001011110100110011110010011111001001111100100100011011011011011100011110111101011000000000100101001000001111100111110011111000111110000001111100000011110111110001001100100110010011010010001001000100100010000111000011111000011111011010010101110000001011101010101101010110101010011111001011111110010111111100110000111010011111010011111010011001111000110111100011011110001100001000010000100000111110010101111100101011111001011000100101001011100000000010000001000010000100000010010100101001000111000111000111000011000000110000001100000000111101110011111011100111110110111001110011111110011111110100000011011110111011110111011110100110110101110110101110110100101100100000001101010110011000101100110001111110010010100100011111011011111001110111100111000111001010110010011110100100010010001000010100010100111010010110010011001100001110000001101101010101010011111100010110001011111101100000110000001001000110000110001111100101010110001101011101111110111011010011101001110100110011101010111101010111101011000100110010011001001100001011011110110111101101100001010101010101011000110010001100100011001000001110001111110001111110010000011110100111111010011111000101001111100001111111000011111111011100001101100011101100011101100000011001101110011011100110100111010110111010110110001000011011111111011111111011111100000000001110011011110011011110011100011111110010011111110010011111110010000110001101100011011000111001000011100001110000110010000111000011100001100110010101100101011001001001110001101110001101110001110011101001011101001011101001000111110000111111100001111111101110000110011111100111111001111001110101101110101101100010000111000000111000000111000000001011100010111000101101110011101001111101001111101010000101110011011100110111001000110010110010110101101011101111010110000100101010010101001010001110100101110100101110100110001010101010101010100101101101011011010110101000100001000010100000100101001010010001100001100001111100001101001101001101100111010111111010111111010111001111001010111100101011111011101001111011111111110111111111101111100011110110001111101100011111011000000011111101111110111111000111000111000111000011101010111101010111101010100111000101111000101111000110001110110100111011010011101101000010111000101110001011011100100110010011001001100000110100110100110100011010101110101011101010100011001011001011001001000110100011010001100010000011000001100000000100111110011111001000000110100110100110100001101001101001101000011011011011011010101100110100100100001101100110001011001100011111100100101001000110011001001001110100000011111110100111110100011111101010100101111011000001101101110010111101100000010111000001110010101001001111010110001001100100110010111111001110101010101001110011100011101001011010000111001010001101111111011110111100010011110101000111100011000100101001010010010000111000011100001100111111011101111111011101111110000110011011000111011000111011000100110001101100011011000110001111111010001111111010001111100011000111010011111010011111010100001111100110111111001101111110011010011111101101111111101101111111111001011010111101001110001100101000101000101000010011011001101100110100111110010011111100100111111001001001100010111000101110001100011101101001110110100111000010001111100000011111000000111110000000010111100101111001011101100110011011100110111001101001111001100111100110011111100010001101110111101110111101110110010001001000100100010010101111010011110011001110111110001101011101100110101111000111011111100000111101010001010010111111001001010010100100110110110110110110110110101001111110111101111110111101111110111100010000111000011100001000011100011100010010000000100100100010110001011000101001110011011110011011110011010011010101110101011101010100111111111011111111111101111111100010000110010111100101111001011001111110100011111110100011111011110000100001110000111000011101011111110101100100100101001010010011101110001110111000111011100000110111001110111001110111001001001110100111010011100011111111011011111111101101111111100011001110101111110101111110110000011110111100111101111001111110100000011110000101111000010111100001000010100010100010000010001111000111100011100110000011100000111000001110101110101001110011011011001000000011010101100110001011001100011111110111100011000010010100101001001111100111111100100011110010100011001101100100111010010001011101110101011011010000100110010011011001101001110110111110110101110111101001110011011100011111101010100111011110010001011000111001111110001011000101111110110000011011001110110110110111001001000011011000100011011110101000111100011010101000101000101000010010001001000101101000010111000101110001011100000101110001011100010111000001010001101000110100100011111110001011111110001011111111010110011100111011100111011100111000110100001101000011010000000000110101100000000110101100011111000111110001110011101001111101001111101010000100010010001001000100001111011111011110111110111101111010011011111011011111011011110100100110110011011001101001101100001101100001101100000010111101101111011011110100010110010110111111111111101111110100110101101000010000100000100101110010111001100001110001101110001101110001101010111001110011110101101111111101111111101111100001111110111111011111110101110000001111101010011101001110100110011111010011111110100111111101010000110010111100101111001011001111011110111110111101111101111011010111111101011001001110110011011000110011000001011100110111001101110010010000001000000100000000010110010110010111000000000010001101000110100010100101110001011100010110111101011111111110110001000100100010010001001111111011010111111011110001110110010000000110101011001100010110011000111111101110001010001110100111100111011000101001111101000011100100011110010100010111101011000101101100011001111110010001101000000111111011010111101110011111100000000111011010111100000011011111000111111110000011111000110111111110011100110100001101001101011000000101001100100100111001000110011001111001110001110111110110000111111011001111110101101000001001111010101111111101010101111101011111010111110001000000100000010000000010100101010010101001100100111010011101001110110101110100110101000101001011100101110011000010101011010101101010100101101001011010010110100001011110110111101101111010010011001001100100110000111111110110011111111011001111111101101001100110111001101110011010001010001010001010100100010110001011000100001111100001011111000010111110000101101011100010001101011111111110110010010001100101111001011110010110011111111101011111111110101111111111011000000000000101110101110101110011111101111011111101111011111101110100101111101011111010111110101011111111100111110000101100001011000001000000010000011100011011100011011100011100110011011100110111001110000110010110010110011111111111011011111110111100011101100100000001101010110011000101100110001111111011100000100010101010110100110010011111000111111101000111111010110001010011101010010101010001111101001100010100001100001110111101110000010011110001111110111011111100000100101101011000111100100000111101101111110000101111000011001111100101011110100111111101100000101110001011010010111010001111010000110001111111111010100011011100110111001111000001001011100010000111011110011110101011010011110011100101011111111010101100100011001000110010000010100011010001101000100100100010010001001000001000101100010110001010010110001101100111110110100100010010001001000000111110011111001111100010011101001110100110100110010101100101011001010001101101101101101101101101100010000101000010100001100010110010110010110001100011011000110110001110010001001000100100010000101010010101001010100111101011001100110010010100100011101100111010110010000101111010001011110110111101101111010011110001001111000100111101011110001100001100001100000010100010100010100001101101001101101001101011110010011100011111011010111011010111011010100111101101011111011010111110110100001111100011011111000110111110001110011100011111100011111100011110101111011100110110011111111111011100110001011001010111000011010101100110001011001100011111110111000001000111000101110001011110011100011111110101011101000011110100000010111010010110101101010010010101101010110011000011111101001111110001011111011100000101101101000111101101000001000000100000111101110111110110110111101100010010111110100100010111100001100111111010011010110001001100101001110011100011110100101100100011111011110000111000100111010111111101000110111011011011011011011001101000111010001110100010011001010110010101100101000111100110011110011001111110001000111110011011111100110111110010010001100101100101100100111000001111000001111000000001011101010111010101110101010111100110111110100111000111000111000011011000011011000011000010001101110101101110101101110100010011111001111101000000111110010001111100100011111001001001110101011110101011110101100011111101000111111101000111110111100001111000111111100011111110001110001100001100001100011111100011011111010111001011001011001011001001100111011001110110011100011001011110010111100110000110010101100101011001010001010001101000110100011010111101001101011101000111100011110001110011101110001110111000111011100000111011110011101111001110111011001110111001111011100111101110000001011001011001010100101000110100011010001110101110001110101010101101101001101101001101101000011111101111111111101111111111101111000111101101101111011011011110110101111111101101011001111100010101011001100110000110101011001100010110011000111111101111000010001001111101001110100010011111110011011110011101111101001000100000001000011000001001100110011101001100001101101001100001110111001001010011100010011000101001111101010011101000111000111101011100111111111100111011111011011110110110111001001011101000110011100001101100010000011110100101100100111111011111001101111011011110011101101110011011000010110100110110101101011110011010111100101000010100001010000001111111101110111111110111011111111111111100010100010100010100001001110100111010011100001101001101001101000110111100110111100110111011001111011101011110111010111101110101010111101110101001110101011000000001101010001001000100100010000111101111111111011111111110111110001101010111010101110101000011100110111100110111100111000111010111111010111111111100000001000100100010010001010010011101001110100111000101010010101001010100001101100101101100101100001100100010110001011101011000100101110111011101111110011010010001000010000100000110100001101000011010000001111111000001111111000001111111100111000101000101000111010101101000010101111110100111111110100111111100000100010100010100010100000100001000010000011000100110001001100010000111111110011011111111001101111110111000001010001010001010010101110011110100101011111000010111110000101111110110011111010100000111100101110101101011011010110110101001111110101101111110101101111110101010010111110101111101011110100111110010101111100101011111001100110101110100110010110100100101001010011011000011111000101100100000001101010110011000101100110001111110010001110100011111100000111010100111000101001110010001100011111101000100110000100101011011101000110011011001111110100000011011100111101111011101101000011100100111001000111000110000110100110110110101010111101000100111100101010101000101100001000010000000010010111000101110001001010010111000011100111011001010111001100001101100001011010011011010100100000010000001000000001101110111101110111101110100010011101001110100111000010010100100000100001000000010001011000101100010100110111010110111010110111010001110111110111011111011101111010010111100101111001011110000011010011010011010001100000111000001110000010011011101011011101011011101000101111011011110110111101000000000011011101111011101111011101000111111110100011111111010001111111101000001111001100111100110011110011000011101010011101010011101010000101000010100001010000001101100011101100011101100010011011101011011101011011100100111011111011101111101110111101001011101110111011101110110010111111101111111011111010101111111000110010001011000101100011000110111101110111101110111100001010100101010010101001101011100000001001001000001100000110000100001100001100001100000110111110110111110110111110000111000111000110111101011101111110011001111100111110010111000111111011111110000000011011000011011000011000010001110110101111011010111100001100110110011110110011110110011101011100111101000110011111101111110111111001111001000111100100011110010000010111101101111011011111000011011011011011011110101100000000101000101100101100011011010011011010011011010000011000011000011000001011010010110100101101001111111011100111111101111010110100010110010111111000011010101100110001011001100011111110110111010001111101001011100100111111011110001111100010111111011110111110011110011010001111010101110100010011010100100101110010100011000000101110101011101000010100010100001011000100111000010111111101010001001101001010011110010001110111101111101011100011111111001011111011100111111101001100010100010000100000101000110100011010010110101110111111010011010110010110010110000110000110000110001101011100011101011001010100111010011101001100011001011001011001000111110011111001111101101011101010011011111001110001110001110000101010110101011010101000110100110100110101111010100011110001110101100011111000110001010101010101010100101001110100111010011111101010001111010110100101011011110011101011110101101000111001111010101011010111010010000101101001101001101000010101010101010101000111110011111001111101111010100011111111011010001110001110001110010101110101011110101111010110010100011110111011100011100011100000110000110000110000001011101011101011110110010000000110101011001100010110011000111111001001001010001010001101010110100100011100100011101011011101000100111010000111010110111010110000110110111000110110111011010010000011001110101000101101011111110101010110000101110101010101100011110000001110110100111000100001101101101100000111011000110110011111011001111010110010000000110101011001100010110011000101100110001111110011010101100010110011011101001000011011001100010110011000101100110001011001000000011010101100110001011001100010110011000101100110001011001000000011010101100110001011001100010110011000101100100000001101010110011000101100110001011001100010110011000101100100000001101010110011000101100110001011001100010110011000101100100000001101010110011000101100110001011001100010110010000000110101011001100010110011000101100110001011001100010110010000000110101011001100010110011000101100110001011001100010110010000000110101011001100010110011000101100110001011001000000011010101100110001011001100011111100110111001000011001011010011001001001011100111010010101111111011110100011110000111001010110011000111111101110111010001011001011101101011000010110011000111111001100110110001010100101010110101000011010010110100111101000000111010110111010111111010011001110001101110010111110010100011010001110101001101000100111111010100111101111011111110100110011011101111011011111011110110110011111011001110010110010000000110101011001100010110011000111111101111111110001010010101001110100100011001011110011101100110000111010001111010110111010001001110010101110010111110010110011000100111010010111010100001101000011001111110101000010100110110010110110001000010010100100101001010011001111111110100001111110111111111110111011111111111100000110110000110000001100001110110011111011001101011111100101000011000101100111000011111100111011001100011111100101010111000010010100101001001001110101000010011100011001001110010111100100000111010001111010101111010100001110011001110011011110100000011101010011101001111101010000110101001101010010010010010100101010011101010100011011011010010010001101101110000000100100010010001010001010000000101000101100000111100001111110000011110111010001111110111101111110110101111110111000010110111101101011011011110110011111011000000110110010000000110101011001100010110011000111111111101011011000011100010010111000010010111001101100110000110010001100101011000111001110010011110011011110001110011100110111100110011100111000111010110111010110110001100010010101001010100111000011001101010100000100101110000000110100110110110110001100101110001101000010010000000101000100001000000001111011010111101101010010100010100010100001000011100000001011100111101111001111110100001111001000001111111100001111111010010111111110001000100000001111111000000110101101111001111010111000111000001101101101101101110101110111111101110010011100010010100100011111011111110111000110111111001110010101100110001011001101001001000011011001100011111100111000001000011010011011011010001001010100110010010100011101011111000111111010111001110010011110010111110010010011100110111100110011101001000110001011110110001100100100100101110010111001100000110010110010110110001101101101101110000011100011100011011000111000100101111001100101010011100100101110110011010101010000100001000000111000100001000000101000100001110110111111101001001001010100000010100111010010011001001111101000111111010100111110101010010110101101101111001000001111011101111110010001111011110000010101010100010110001010101011001011001000111000111000111000111100111010111111001010100000110010110110110110001000000110110001001011110011000100010111010110011000101100100000001101010110011000101100110001111110001101100001100101101001100100110100001101001111010000001100010011101100011000100001110010011110010011110010010011100101111101000011100111000110001101100010111001011001010011101000010100100010101001010100011101000001110100011011011110011011010111110101101101110001110000010010111000111001101011100110011110011110010010100001000000100001000010100000101000101000100000000100001001011101011000010101111001001010010010101010111000111000010011011001011011100001111100011011111110100111111001010000101110101110101100011110110010111100001111110001110001010000011111000011100010010101000000011110000000101110010100010101010000001000010100010110001101001110010101101010000110100111001001110100000011011001111000010110110011001000011100000110001001011001111000001010010110010000000110101011001100010110011000110101101000101001110101011010011001100110011001101110011000011101001111101011011101010100111000101111001100111001000001110100011110100001110100000011001110110010011101001100101000110011111010010001010101011001011010101100001001100000101001001000110110111000110100001001000110110000000111100000001011000111000111011111101111101110001101001101100000100001000000101000101010101010001000000110010001001010100010000001001010100010110000101000101000101000001110001000000001110001001010010001001000101000011010010110100001010000001111100010011111110010111111110100000011111010000011000010001110111111111000100111101100000001000010010000011011010010110100001100110101001010011001010010110100101100110100101000011101011011100110000110011101110101001100010000111001110110011111100101000101001011110111110111101111100011100000111100000011101111010001100001011110110011001101101101010110010000000110101011001100011111100111010111000010010100101001001100101011001101110011000011110100111110010011110001100011100101011100101011100100100111010000111001111111010011001100111011001111100100100101000110100111010011000111000110100110010001001011100000001001010010100001110110100100110110000111100101110001010100100001000000100100011101011111100100011101000010000001110100000010011001110001110000011011011100011101100110100010100100001001000001101101110001101000010000100001110000011100010100000001010001000010010111101001101101101001110111111101111101001000101000000000100000110100001100110110011000011111111101001111100010011111110010100100000110000101000111000110101001111011011001110010011110011111110001110011011100011000011110110000001011110011100100011110100010010000001110101011110011110010110111010010100000111011101101111100101010010011101110100001110011000011001001101110101100001000110110001101111011100001111111111110010101101100110101001110110011000101100100000001101010110011000111111001100010010000110110110110110110011110011101111010001111000111001111111110110111111111100011111000101001001100110101011010000000110100110100110100001101001001011011000110110110110110100001110001001011011000000010010001000000101010111011101010111000101000011100101011111011001101110100010010001001011110110100100000100000110110001101101110001001000111000110110111000000010010111011101000101000010101110110100101100001010010000010000111000001010001001010010001001010000101000001000010100011110111100110010010100010000001001011100011100000110100110100110100001010001010101010000110100001100100010010010011111111100111111111110001111110001000010000000111110011000001010011101000110100000010111111100000110001110010011001100011011001010001000110011100011001000001010001010100100000001000010110001001010110011101101001100111001110111010010111010001000110010110101010101001101101011100001011011011100010110010101101100111101001011100111111101111100010001011001010100101110111101100110001111111011110101100110011010100111000111000111000010100101010010101001101110111010110000101010110111000110111101000111000110110100000101010001100101101100011001011001011010000110100110110111000111101011100111011100111000001101001101101101000011011011110111110101100010010111011011100101000010110110111101001100010101001101101110001110100011011001010101101111100001110001110001001011101111110000111101111001111110110110111000100101110100100000001111001101011010100111001001011101111111011101011100000101100101000100000010101010000101010011001110110010001101000100110100011101001111010101001101110111110110100110111011000001011101100000111001011100101001101100111001011100101101000001110100001001100011011001110100111010101000011101100010011011010100001100010011101010011001001001111100010111111110100011111110011000110001011100100011000100000100101110010110011011001110101111011001100110000110101011001100011111100111011100000000110100110100110100110100010100011010010101001000011011011011011010001110000101110000001110000000010010011101010010011110011100010111100100011100011000011011010010111000111101101101110001001101110000011101001101000101110101000111010010001110011100000111011111110011001110010101100000001111000100110101111101000100000010100011110101110101000001101011000100111110111010000111101010010111000101000011110110100100010001010100001010001010000010110010101010101000101110101100101010010000110111111011111000101110111011011110001110001100110101010110010001001010000101110011010010100101110100010010011001101001110011100011100100011100010111100100100100011111101111011000001001101001110001011011100000111010101110001111001111000101110110100110100011000010101101011011010100110111010110111100111000011001000001011100010101001000010011000010010010100111010011101000100011010011011011010000101100100001011011110101100111010110111110111101100110001011001000000011010101100110001111110010100000100010100001010011101000000100111110011111001110001011011010010001011011110101111101110101010111011111100011100000000110100110110110110110110010100101010010101001000011011011010011100000101110111111010101001110111101111011110111101101000011010010110011111100110100111010100110010001100011000000100001110000010000001110100000001001001101101110001110001111011010101110111110010010001001001010110001111100110100000000100101000000111000111000111010000000100100111011101001001111100101000101011111011000011011010011101000000011010010010001010101010101000001000001011111001100000100011010000111000001001000010100001001100000100000101100010000000010010101001110100110000011000011000010110001010001101000110100110010111011101110001000111001010000101001010101010010011011001111101010100110010101110101111101000000111101001001100011100100100101101111000111100011000010110110110010101111000011011100011011000111011001000110000111101110101101100100001010110001000110000010011111100110011001111001110101111100011111000110001011010110110111100100000110110011110110000110110111000101000101000101001011000000000110100110110011000101100100000001101010110011000111111001010100010011010010010101000010100011010000001100100011001101110010100011100110111100110111100110000111001000111001011111001011001100111011010011110011110011111101101011111111000011111110110000011101110001110000101110001001111111011000100000000110101010011101001110100110010101000110011010100001010011101001010100000010000101000011011111000111011111111110000111110111010001101000011111010000110100110011010101100101110010110001010101000011101010000010111001000100110101111010001010111001110100001010001001000010000111010000010100100100001110100000001101001110101000011000010101110111111000000100001000000101100101000100100100000001011101010100100010010000111000010000101010101010101010010110101100000001100000101111011011010110110100001100011111010100110100100001011001010001110000101001010100011010101001110101101100011011010000000110000101010000111000010110111101110110001001110111110111011100011100001100111110001101111001001111111101010001001001100110110100110011101011011101001111000101001000110111000011110111011001110110100111011110011100010000100110010100101010000001111101001111111100000111100110000110100101101000011010010000100001111010100101101001111011100011101101011110111000001010001101001010100110001011001011001011111010110111111101100110110011000101100100000001101010110011000111111001001110100000100101010011011001110100110100110001011100100111000110001110010111110100001110011000011100101011100101011100110000111010100111010100110001010010011001101010110011010001101101101001001000100001011101000001111100010111111110011111111110010100101111101011100110111100001100000110111111110000101111111010110100111000011010011001011001011001001010101101010010100100001100101100110101000010011011001111100100100101110001011110010001110011101101111110110110111011010000111100101111111100000111100111000101010101100110100111010111101001001011100000010000001001010010110110111010001111010100001000001010110001101111101110101000101010101000001000000100100010111010101000001111100101110101100001010001000010010011000001101110011011010000100100010001001000010001001001100110110011000001010101010001010100110011111101010011010101001100111110010111101010100010111011111001011100111011100011101101111101111100010111011101101111001010001111110001011100011011100111000100000010000010101110011010011110100111001111001110111000111011011110001000011111000001111101110011111010111100111111111100011111001011111110101110010100011010101101010100111010010111010010110001000011000101110001111100110100101001010100110110100001000011100011101001001000111111000011100000101010100111101110001111000111111100010000111000000110111011111000000000110110111000000101000110100101010011001000101100010010000111011001111001000010001011001000000011010101100110001111110010010110100001110001001011100001001100100110110011000011000110110010011100011000111001000111001100111001000001110011101110010111110011000011101000111101001111001001001101010010010111001010000110110110100111000001001011100010010001000101011010110111110111001101000001110010001110010011110011110011111000101111110010001111111001100011111101110111111000010111110000110010001101000100100011011110101010111110011100110101111010011000111001001010010001101101100101100100101000110100111010000001101000011010001110100100011001111110100011001010001000010100010010001110011000001110000101100001000110001101110110001110101011101011100101010110101110101000100001000000111000111100101100000001010100001010000000101000001000000111110011111001000001011011110010001000011001000100011111101011000010110010111010110001001111100111110100100010010111001101100111000100111110011111001111000111111011000010101001100001111011000110111010001010011101010010100110011010011100100110011110010011001001110101001100110100101101010011010000001111110100001111011100011110001010001000010010110110011000111110011011100110100101010101101001100100111101000111100100011101000100111100010111110000101110111010001111011011111110001001110111101001111101010011111011111111101000000010111011000010000010110111100010110000000001001100001110000000011010010110101011001110001010101011001101010000010101010100010110001100001111011010111000011000110001000000010100001010100101010110100110010000000111111100000000101001110100111010011001000001100000110000011011001111001000001001011001000000011010101100110001111110010010000000001001010100101010011001001010001100010111001000111011000001110010011110010101110010010011100011111100100111101000000110001001100010011101011100100111010011001001101000110010110010111000001101101110001000000110110100101111001011011000101001001011101001110001100100100101001011101100110110000100110110110110100000111110110101111101110011111011111001101100011100001011011000100111101111111111011101011110111110000101110101101111010100111001100100111100110110110110110110010011101001111100111100010010100000000110100110100101010011101001011101001011101011100011100011011011011000110100100101011000010000101100111111001011100110111100101110010010011001001011110101000011010101110100111101001100010010001111001001010101000001000010010001011001010000000111111011111001010100100000101111110111110001011100110110111100100000100101010011011001100001011011010010001000011000100101101001100100101010101100110100100010000000111111010100001101000111010100100101000000111000000010110010100011100001111000101111101011111110111010001110000001101111001101110110011111110011111111000110111110101010010010001011010010000100011000111110011001101000000111111000101110001011111010001001111011011111110110100111101011100011111110011011111000110111100100100100010110000100110000010110101101101011011110100110101001001010101010000111100100011110110110111101101000011101100011001011110100000011101000011000100111010010001110111101111011100111101101000011101110111110111001111101100010011110011011111010000111001110000100001000010100000101010101000110010010100011001111101000100010101010100010000000010010110010001011001011001010000010100010000100000101010110101001010101000101110111110010111101100110100101100001111111111101100001000101100111000011111100111011001100011010111100000100010001110001101100110100111101010111010011001110110001100011111101011100111000111111001010111000110001110010001110011001110011100011000101111011000110010110010100001001110101001100011011101010001110000011010010010111010110110010110100011100011110101110010101110011011010011010110101110100011110101011101000111000101001110110011001110010010000000010111010101010110001011110110111011101101010011111110000011111110000011111111111000001111000000111011110011110000011010111000001001010101000110100101010010001010000101000110100010010011001001100100110100100111110100011010011001010101101010010101010010010011001010101000100111110111101111001011111100101100111010111111010111111010011011101111100101100010110010110000101110110000110000010100011001011100101100110001111110110001110110000001100101110001101100011111001011101010000100001001111110101110000010010110100011101101001101111101101101110010011101001110101000000100101010011001001101001101001010010101001100001001111101001010100100001101101101001101000101111011011100010001110011110111011111100011111110101111001111110000111110011101110011000011100011011100101011100111100101110011011011110110100001101100101101100001011110100111111010001111101110011111000110001110101101110100111100011000111110100111111101010011111011011001001111011011011100001000100100010110000110011111000010111111110000111110111101001001000100001110111001000111111100010010000010010101000111000110000010100111001110101000100101101111011100001100000111001001111001011110001100011101000011101010111101100000111000000111000001110000110011110110010111101100001111000101001010001101000001001001000010100010010001100010100011001111101001100111010010111010101111001100000111110011111001101100110110000110110000110110010001011111010111111110000100010011101010000101000100111010100110001001110100110010101001010101100111100111011110011100010011101111100010000010111111101100110011011011010101100110011000011010101100110001111111111010010110000110100110110110100011010000110100001100111000111010101111011000111010101001110010011110011011110010110011100100111100111111100111100110010111100010111001100001010001100111110100010010101000110010100100011011010010100000010010111000100100010010111000110110001110001001011101110000001000001101000010011010110110001000111010001110010101100010000100101010101100001111010100111010111011100010000010100010000001101101001010100001101000111001111100110000111111111011111111000100111110001010010010001000110100011100110110000110000101101100110010011011001111101000000101000110100111010101001010100101001110100110010101010110010110010010101001010011101010100110100101101010011010011001100101111001100110011010010111010101110101011011000110001101100010101010000110101001101001111010001000111111100010110001100001110110010000110100011100001011011110110100100001100110110010110000011011110100110011011101000011010000001001000100010010000110011101011111001010110010100011100011011100110011101000100010000001001001101101001101100001011111000110110000101111111011101100111100110111100100011100110100100110110100111010001001101001011010101000011010000110100111101000100111111010111111101111111111011010100010100010010111000011001010110011111101000000111001110111010001111010110000110100011111010011001111110101101111100000011111101000100110101001101010010011000010111000101111011011111000101101001011010110111100000110000110000111110001000101101101000111111001010101101000111001111001100000110111111110111100001100011011000110011001000101000100001010000111100010111110010001111000110001101111101100110010010010011101011111101011011100101000100100110010111101010000101010010101010110010010001101011010110000100010111111110000011011100000011100010100110111010001100110111001111110001110011010011100100111010101001111001111111101001111110100000011000100110001101100100100110001011100100011001101001001001100110011001110001001100100110010011010011110110110111101100111111011011000010110010110101100101110000111100001111111111010101010000101011111111000011111111000011111111000011111111000011011001111101101100001111110011111110100010101010110011010100001100110011001111110011000011100010111100011111110100010011111010010111110101011111101000100111111101001111110010001111100101100111110100111111101010011111011011001110010111110010001110100110011001110110011001101001100101010010100010110100001101001101000000110100111000111010100011110110010111000110110110110001101101111011111001110101101010010111111001001001010110100110010110101101011011111011110011101000000111010011101111110011011101001011001001110100000110101011101001010010010011001000110011011100010100110110101110110101110111000000100101110001011000101001010100011010101001010101101010101110000011001011010010010010100111010010101010100110001111100011011001000001101010111010001100101000000111000100100110110100110110101110111000001101000111010010110100110001010001011001010000010110010110010110001010101101001010100100010100111010001100111000100000001100001011100101000110100101010001001000001011111101011100011010101010101001001001011100110010011110010011101001111101000100011000011111001111100011110111111111101110101111001000001000100011111101100000110001111100100111001011001011010110001011000111001100010111101100011001010001011110010111101101101110011011110011011100011011100000111010110111010010111010111001101110011101100111101110000010111001101110011011111100110110001110110011110110001001110110111111011011011101101100010010001001000011000001100001111011010011011010100010110010101011111000100111011010010110010100010000110100110011000010000111000110100001100101111011100001011011101000100101110011001001001001011101011000000110000010010111111110000001011111000011111001010010000010011101100011101100011101011100101110001011100110111000000110010100101001001110100111100010011101011000111101001011100011011110100000011111011101111100110011110011000011111001010111110011001111101000100110001011100011011000101001101010110010011001010001100111111001111110100010001100110100011010011001100100011000110110001000010010001011010010001100011000011110110001110110100101100110100111100001101100110011000011010101100110001111111011011001000010010100101001001010100011001101010000110011101101000011001110001110100001110100111110100010011100100011100010111100011100111001101111010000111001111001101000011001110100100100101000110100010110010001101001101110101101010100010111001110101010100100011101001010010111001010111101001000100011010110011111000001011101001000100101110110011001011010011110101001000000011101011011000111111101000111010011111101001010101100011111110101010101101001100101101001110101011011100101001100100011100010100010101001110001101110001011110011110011111000111101101111111100011100111101111011111011101111111101001000010000111000101110001110001110001000000111000111000111011011100001111101011100110111010101110110011000001110000001100001000010101010101010100000100001010001010000101000010100001001111001110001101110010101110001010111100000001010010100100100110010011011001110001001010100101110010100001011001010101001001110110110111000010110111001001111000000111011100110111110001111100100011111001101111110101010011010001101010010100110001111110111111100000100111100110111100010111110100110011110110100111100010011110000000011010000110011011101001100111000111111001100111010001001000000011000100000100111101001011100011111101001100111110000101111110110011111110101000011111000010111111011010101110010010001101000111100011100100001010001011011100000110101001101010011001101001110011111110001011111101111100100001001010010100110001001011001101001000101110101101100011110000010001011001011001110000101111111011111111000001001000100100011110110111001001111100110110011100010011001001100100110000110011101101001011001111001011111110111101010111001000000100011101011100010000101110111110001111101111111110011101111001110001110010101110011001110010110010101001010100011101000001111011110100001101000010010010011010011110100101001100001101010111010011110101010010101001010101101010000011100011100010010010110111101101101001000001101001111010011100110000111110001011111111010011111111001110010001011011010010010000011101110011110110100111011101110110011110010010111010110010000000110101011001100011111111110011011000100110010011011001101001111100011011110010011111100101000111110111011111101111111111011111001101010011001111110101000010100111001111101010100011010011010011100000110110100101001000100101110000000111000001110010101100011010000101000010010001110100111111001010000111000000011100000110111101011011000110000101000100011010110001001010101110001001011101000001111010000100010101111001000010101001111010101010100001011101111110100001001010100010000001110001001010000011010110100100010110000101000011110011001111110000111110011110011101110001110110110111011110000110110101110000111101110110001110001110001100100010000110110000010100010000101000010110110101101011011010000011011011100011101110011011100000101001010010111000011011110011011111011011110000110100001101010110010010011001001110010011110110000001110001001000001100101101001101000101001010100011010001000100101001101010100110101001001011100111000111101100111111010111111011100100111111010010010101000011111110011111111001011111110100100011001011110010111100110000110001011100011111000101001011011010110101101101010011110110111111101101111111001000001100001011000010110000010011100001011101101011110001000001000010100010110001010011101001010101010011001110110100101100111000111010101111010111111010011001101101111101110101110000010010110101100100010110101000111111110110100110111100001011010010000010110000010001101011111011011001100101010101001010111000111000001010000011111110001111011101000110100001100101011101000000100101111001111111010110000101010100010000010011101001111101000011101000000111110011101111101000111111010011001101001011010011110100010010100101010001011001001110110001110101111100011000110100101101001011010011001000110100100010001100010011011001100100110000101010110101010110110001011001011001100000000100101010100100000010000011000011001000000100000101111100010110101101101111011011000100010110000011000001001001001110100111101010100111111100100111111111001111111111100110010010001111111000001001000001101110011101101011101110111011001111001000111101011001101001001000011111110011111011100001110001110001101100011011011011011011000100001000111111101100110010100001101011101011000000000110010011111010000101000000111001011111001100111010101001110001011111010011111000111001010011100111110101000001101101110001001000110100111000110100001101001101101101001111011001111111011100110110001110001111010111000111111001110101100010011011100111011100110101011110101011111000100011101000100110101110001000110101010111001111101010100111101001110011101010101111111111011010010000001111000000000011000011101011101101001000001000011110011000111001111001010001000010000001010101010101010000010110000000110111000110110111110110111001101100011100001011011001010101110111010011010000011101000001111110011101111100010110100001111011110001101010110010101010110001011011110110110101110010011001111110011101100111100110100101101001111010000001000011010111011011001011111010111001101101000000010010100100100101110011101001011001010011011011011001001110111011111000100111011011100110100101101000011010100000111111011000011111100111100001111110000011111000011001011110010110111101111000011011101111100000011011110000010100010011010010000110110111001001111001011010010110110101110100010100011001110100111100100011110110100100100000011100010001000001001100000111000000110000110010001101000100100010100000101110101100011000000110111001111011011000100101110010011101000100110100111100110011101010000011100010000101000001010001111100111111001111010011111101001011110011010011100011111100100111100100100111000111111010001110010010011111010111111110110011111001011001110011101110100001110101010001100101101101001001101000111010000110100000010011111001110101000100101010010101011010100001010010101000110100110001101101101100000111111011111101111110010001101000110100011000101110001011011110110110011101111101111111100001110000100100010001111000110001001111100111010011100010010111001101101000100110100001101000011010100001100110111010000110001110011100000111011111011100000000100010111110101100001001001011100010110011000101100110011000011010111111001100110110100101001110011010011010011010001001111101000010011100010011101001111100101000100110110010111001011000101010100001010100101110011011101110111110001000111100011110110100011110110001110001010011111100011111111000111101101101101101110100000100111011011111111011110111011110000111010010111010010110001000011100011011110100111111010000000100101001011100011110101001100011100000011100010010110100111100010000001011101001000101000100001010001110110011011011010010011010110101001101111100010110000000000010010110101100011101110101001010000010001101011100111010110010000011101010111011100111110101101111110111000111000100101110100000011110010000111000000011111000010110010101010000010111101101111111011110100100000110000001000000001011110110111001110000000001010001000010100000101010101100111010111011110010000010100010100010000001101101000010100011110101001100001010101100001101101110001110111000010011100111011100110111000101101000011101101111110110101111011100000110010011100010111000110001101000110011011010010001101010011010100100101100010100010101010010001100010100110110100011001000111011000110011110010101001110111110010000011111111000111111110110001111111100011001110101001110101011110100100010111110110000011011111000011111001011110001000011000100111010010111010100001100110111101100011000101001011101110111001101101110001010010110110101010000100000110000111000100000111110011111101100000110111110111011010011101111100001100110101001010001001101001011001110110001110001000010100010100000110011010101101010000111101001011110010111111101111000110010101100101111101001100101000001010110010000011101010111000111111111101001001010011011011011100001000000100001110001000010100111001110100110100100111110100011010101001001100100111110011000010010101110101001001011000110101010001101001100011000011000011111100100000010000111000010000111110011111101111110001101000010010010110110100011110001000010110111101101111011011000011010101010101101100110101001001001110100110010011011001111100111000100110110011011010000000110011010001101001100011000100001110000010010001111000111100011000110010001100100011001011001110011111110101001110011000010111110101111001011111111010111010100101010011101100110001011001000000011010111111001100000110011010001010011100000110010110100110010010011111001111100110100100110110011001001001001101010111010101110101000010011101001110100101100101010010100111010100000100101110001001001000000011111101111110001000010000101000001011101011101111100010001001000100100010111111110101111111100111010011001011001001010101101010010101000001010001000011001001110111100111011110011101101110011001010110010101100100000110010011100100111000111101011111000101011101000100110101101001000110001000010000111010011101110101001111010011001111100101100010000010110100111011100010000100011010011010110001010011010100001110001111001110011011110010100001000010000001010101010001010001110111000000110011000100100000100101001011011001000000011000010111001011100110110110101101000010010111001011100111100110111001110110011101111000010011101001111101000000100101010010101101001000011011011001100010000100000110000101000000000101000101010101010001010101001010101000101000101000101010001001010101010010001011001011100101011111111110110100100001111000000000000100000000111011010011100000111011110000011001101000111110111001001111101001011111010010111100100100000100001101000110000111100001010111011001110110111111000010110110101001101100111100001111011010100100000110000111000101001100100111001010110001100011001111110011111100111000101001010100111010010001100001111011010111011101000011000100001110001000011101101011110111111111101100100010111011101110011011110100100000110001111000110001110011001110010001111010011000111110100000010000100001001011100010010011100011111110011001111101011000011010011010101001100110101001010001010000011111010111111100101011111011101001110110001100010111010000001010100101010001010000100101010011001100100100110010011100100011001111000100001010101010000011100010010110100010011111001110100101100011000011111110000010001010001010001010100010100010101000010000111011010110111001001011010110110110101101010010001101000110100011000011010011100011010001100011111000111110001010011010010110100010110010010010111101010110011010010011011001011100101000010100011000010110000111110011111001100000010110010101010111001011010110110100100100000011000011111110000000001011101011001111100001111110101110101100001011101010101111100001100101100101100100010110010110010110101100100000101101010110010000000110101111110011011110100110010010101010101101010110101000010010101001100100100100100101110010111101010100100110110010111101010100100111010011011001111001010100101001110100110111011100001110111101000111010100000010100011010010101001010101000001010010110110010101001001001110100111101001000000001000001100001011011000111011001000011111110110000110100010010100001110110011111100111001101011010011000010110101010110101011010101000110100110100110010010110101101101101000100001111000000111100000011101111000011110010011111001001110100010010100001010000100111110110000001110110010101101011101111000100110101111011101001111100100100011101000001110010010100011110110001110000110001010001010001000000001001010000000000111000111101100111011011110010010001010101010001010000010000100000001000101011111101111110011011100111011001010111111001100101111001111110011100010111011101101111000111001101010011010011100100100111001000111001110111010100000100001000010101001011110010111011100100000111011100111100001011011110000100100010001011000100000101000101010100000010110010010101010010101100010000011101001110110100101100001010100011110010001110011001010000111101111001111100111011010010001000111110110011111100011011110000010010111000101110011011010100011100010011010011000101010100001100100100111010010011100110000110100001101010011010010001100001110001111011010000010100010101010110001101111101101111101110111000000111111100000110000100010111111110110000110000000011101001011101000011100101000100011110111010101111010001011110001011001000001100010011101010111100101000100110110011011101010000101000101101001101000110011011101001010010100011111100000111000110111010111001001101100111010011110011001000110010111101000000110011011101000011001101001011011110111011101110110010100111010010101010000100111110011101001110000001001010101001010100101000110101000001001000111000001111110111111100001100100010010001001011010000100010010001101000111000110101010101101010100100101110010101101010000010010100101110000100110110011001001011001001100100110110011000001110001100101110000011010011011011011001010010011011101010000010111010111011111100100000110001001000011000111110011111001111100001111100111110011111001110110100111111101010100010101000001001010100000101110111110011000001011101010111001101111010010100111010011101010000011111101111110000010111101100111010011001101000101100100000001101011111100110100001001100100101010100111010100101001000100110110011011001100001001010100100111010100001001100100110110010010010011001001011100101100011011011001011101010110101110010000100100001101010111010101100100100100000010000011000001001000000100000001100000100000110000011000001001101111001101111011110000100011010001110100001100110000011001101001110100100010010111001001110101000011010001100000110000110010111111110000001100000111110101100111000010000111011011000110100100100001011010011010011011001010011101001010101010011011010111011001111011000100111000001110111110110111110001111001110111101000111110100000111101011100101111100111100010010001011101110111000010010111100000101011010111001000000101111001111001100010100100001111010011011110010011100011100011011011101111111101110000010000001011001000010100001000101011111101111110001111110110000101110001111111000001010100001011010110110100100011100111011000110001101100100100110100001101010011010100001001110101000010100010010001111010000101000000101101111000111100001100110010001100111011010000011101110100000010010001001010010100001011110110111100101110000010001000110000110010001011101000011100000101100101110101110111011001101010011001000000001000010100010000001000010100010101000101010111100111011111100000011101111110011011110110110100111011000100001000001110111100111011110111101101010011100011111100011111100010100101010010100001010011001000011100001010110100001000110100100010010000010000001000001100001100101010101101001101000111000010110111111110111110000100001000010110001100111111010001110001110010011101010001100101000100111010100101001100001100111111010010110100110011111011100111100101111111011111001001101100111110100000011101001011101000011000110001010001101001001100100101101001011100110111100000110011010101101010100100111110101001010100000110100111000100000110011011100101111010001001010100101010010101010001010101010001010000100001110000011000101001000101100011110000010001001010010000010100010110010100001011011110111100101110100001010001001000010011011001010011001001010101101010110100110011001011110010011100100000011010011110110100100101010001000101100010110001110010000101000100100001100010110010110010110000101000101100101001010110111101101011100010101010110010110100001000010000100000010110010101010010001011001010101000001000100100001110001000010010001000111101101000001010101010101011000101000110100011010010001000011100001101010011111110101101011101111010100010110011000101100100000001101011111100100010010000010010101010010101001010100010010011011001110100101100110100111101001111010001001001101100110010010110010100011001111100111100011010011001011010011110001000100010111101011001001101000000000000100100110110010110110011110110101001000010100001110000110011000110110001011110101100001101001100110101000011010011110101001100110100101111001011111110111111001110110001110101101110101000010000000101010101000011010100110100101100111100100011110010001011010000100011010001101111010110111100111101011110101011011111001101000010100010100001010101101010010101010010101011010010101001000110110111110110111110110110001110100101110101101110101110011001111110100001100110000101100010011100101011100011110011010101100001101001000100100010000100101000110101110011110010100101001100001011001010100011000010111010101001011100110010001000101001001111101000110101000010111001100100010001100010000001000001011000001100110011010001110011000011010100110101001010100001001100100110110011110010010111001110100111000010000100001110000110111101110110111110000100011110111010111100011011110101111001111111010001111100100111111010010001100011011001111110011110010001111011010110110100001110001111110011111110100100010010001000110100010000110111010111000000100000000011000100001110111010000100001000010100011101000100011010010101011101100110101010100101000100001000000101000101000101010001000010100010100011110100110001011100000000100101001000101110101100100000110111100110111011110111101001100010111000110111011000001101101011101100101101100010010000100111111011111000110011111100111011000111001010100101000110011100001111100101110101010011101011011000100111010111001111110000011110011111111001010001100011111001001110010000010011001111101011111110010100001101001101101010100010010110110111000010100101010011011001001101000111010101100111000101001110100011010001001101001110010111001010001001011100110011010101000110000111110100000000010111010110011000000101110101101000001000111110011000100000100100011010000111000001001011011110110110101101110001100001111100111110001100101011001100110011000010010111001101110101010010100001010101100110000100111110010111001101000000010000010000000111111100000100011000010111011111100100010010001001000110000101110101110110000111010011100110000101000010100101011101101111001100110100101000011101111101000010101000011100011100011101101001000111010000000110110110110110010010110101101101011001000001000000011111110000110001101001101000000100001000011111000101001010100101010100001000010100001010000001011001101001101000011011001000000011010111111001001111110000110110110110110100010011101001111100111000100111010011101001011001101010111010101110101000010011001001010100101000101000110100001010000011110101110110001110110101101010010111101001110101111100101001111101011010101010100110000100100001010000101000110011100011000001110110001110110000001101010011010100110100100011110100111111010010111100111000111010010111010110111010101001110110110111011011111100010000011100000111000010011101001111100110100011111001111101000000001001001110101001101001100100010110001011000101110101110000000001010101011011111010110101100101100101100001010001010001110100111110001010101010010100101010100001100101011001001110011010010010111001001110100110001101101001000011000011110000111101100010011010101100100111010011001010011101001110100100111100011101100101001111000111000011010011110000000111001010101010100010000001111100101010101000001010001010101010000010101010100000011011111011011011111000011001101001111010011110101010001111110101110101010010011101001111100110100111010001110001011110110000001001010010100100101110001011010010001000011110101111111011101111101101100011110100101110010011110100010011100110111101001111101010100011011010000111000011001101110100111101010100011000100000101010100111111010101111101111011111011010100111111111000011111110011011111001101001101001011010010110100010011101000110101010110110010111111101101101011101100110000101100001111010010001000011101101001011101000000100001010101111001111100110101110101001010111110110111011011001010110011101010011000001000101011100101110011111011101100110100100011011010110110100100011100101001101100110111111001100011011001010110001110010000100110101001001001001101110101011101000000101010010011101001011001111101000011111010000111110011010011101011111001001110100100011000110110001011100101000110101011001001100101000110010011100100111000101001000010100010110001000001010101010101010000100101110010111001110000100001000010100011101010011101001000011011000010000111000010100011100100000110000011000011001000110100010010001000001111100111110011000001100110011001110110100100010100101010100101010000100110110011101001110001001010100101011010101011101110101011011110100100001000000110101010011011001001000001100000010000110001111110110000111111000111110011111001110100111110100001110101101110000110100010000111010111100101000001011110110110000001111001010110011111111101101011010110010110010000100010000001001000110110010110111101110011000111000100001010001010100101010101101001101001111011100011010000100100001010001101001000100001110000101011001110001011101110011111110110110010001011001010011010110000111111111101000100011111000101001101001101001101000100110110011011001011001101001011010010110011110011000101110001101110101100011001000110010001110110000011001100110010101100100100100101110010011001001011101001001111001110100111010110010001110011001101100010001100010101011000111111010100100001000010000001101101101001101000011010011001101010000110110000110000111101101000011000101111011000110001010010100011010000101000100100011010000111000101001100011011000110111010111011101001001110111010110000110000001001000000100001010000111000011110101110001110100110100111000111000111000010101001010100101010000100101110010111001011001001001100100110010010010011111001111101000100100111010011111010100001110100001110100101110101100010010111001011100110000100111110100011010000000101110101110101110001101001101001001001001100100101110010111010110000010001110011101101001001001100101010101010010001011000010011111100101111011011011110001100001111110101110100000110110110110110010110000010011010100110101001101010100101001010100111010101001001101100111010100000001111100111110010101000111110010111010110001101010110010101001101001010101101010101101100101001010100011010011001110000111101111111101101100011110110001111101011101110111111001001001110100101101001100100101110011111010000001010101011001011010001110101011110101111100010100111011100011100010011100001000101010010101010100100010100000101110011110111101111101110011111011100000101101011011011111000001000110010111001010100000110001000001100000000100010110001101011011101110100100111011011011110101001010000011010110010010000001000101011000100010011111011101000001101101000010011111010010101000000111010011111010111111010110001111001011111111000101111110000000111110101011111101100111111011001001011010010010001000100001000011011000100000100111100110111110100111110011110011111010010111110110011111001100001101001111010100101000000100110110011111010001001010001101000110011110010101001010100101001100100110010011101001110001001100100111010011110001100101100101101100011111101011101100000100010010001001000101000111110100000010000100000010100010101001011100010110111101110100010000101000011100001000011001011010011010001001110100111110100010010011101001111100111100100101010010111001010001010000101000010100100001011101111100111111001000010100000110000100010000011000001100010000100000001111111000011101011101111110111010101010110111101111011000100001000010101011110100110000110100100001111000111011011110011100101011001110100100000010111010000000111010100001110110100111001101010000101000000111011101011101110011110110110001101101011100001111011100100011001011001011010000110110110110110110111101001100111101001110000010010111000110110001111100111110011111010110011110100010010010110011001100001101011111100100110001000100110010011101001011001100111111010000110011000010010101101010011010011001001111100110110011110001101001100101100101110111101110000111100010000010011011001100100111000011010011010011011001001000101101001000101001010110101111101001110110101101001111000100001111010100111000110001010111111010110000001010111000000111010100100111010101110101010000010000100000101101101011010110010000001001011100011010001101001011010011110100010011010001110011011101000000100000001010101100000100010110001001000110001010001100111110011100011010100110100111101000100010110010110010110000101010101010101100010101001010101101010100100111010011100111011100010111010100101001110100111010100001010101101010001100100101010110101010110100001010001011101111100010111111101111011011111100111101000011000110110010010010100111010011101001000100001010001001000100001011010110110101101101110011010010110100011101000100101010010101001010011000101110101100101000010111001101101011000111000110010110100110100001010101010101101100110110011110000111100000000111010100111010100110001000011001001110011001100101100101000010100011010100001001011100111010101000000010010111000010111110101110101001000001111011101011110110100111100010000111110011101111101000111111011100001110101011110110001100100100011011000000111101001011100110011101010000110000111100001111000011001110111101111011101111101101110011100101111101011011101011100010100101010100000110000010001110011001110110100001001100001111110101111111111100011111111010111001101000011001110110011010010001011000011011111000100010110110101110000100011100101011100011111110100010010000011000100110100000010111100101111011101101011010111011000110011111001000000001111000000110100101010000000100000001001111100111110011010011000101110010011100010100111001000111001010111000111001110100101110100101100010100110010101100111011001111001001111101000010011100011010000110011101100111100010101010100011010001111100001111111101100011111101101000100000110110110110001110001111111000011110010000011001101110011111100110000100101110010111001101000100001010001110000011111110000000111110000101110111110011111100100000001010001011000100001010000001000001001011010110010001011100100010110011111101011100100101110011101001011001001010110011101001001001100101111001110110010010010101001010101101001100101010110101010110010010000101000000100010100100000001111110111111000101110101100101110001111100101110111111011101110101101000001100111101110000110100011101101100010110000110101101001100101111000101100000110011100000001011101111111010000011110101100110101000011100010010001000010101011101011010101110110000010000100100000101000100000010111011111001010100101101111011010110111001000110100110110111010101101001101100111011111001111100110110001001010101010101001010001101001101101000010100010101101001000100000110000001000000101100111101000110100101100110011000011010111111101111110110001010010101001110100100011111011110111111000001111101101000111010010111010000111001101000100101101001110000101001110100101010010001101010111010101100100100011000011000011000000101000101000100000100011110010001011010100110111001110111001110111101001001011100101111010101101011111000111011101001111010100010011111101010101011001100001010110011101011010100001010001000001001000010101011010011101001000101000110011011001001001001010100100110010010001100001111100111110001011100110111011101110100010110100101101111011011100010100010101010101000111000110110110110001000010000000011011011100010010010011001010000101001000100101010010111001101001001111100111110100100010100111010011011010001010101101010101101100100110010011101001100001100011011001011110010010011101010011101010011000100000110101010101011010000110010110100110110010100101010011101000000011111110000001000000000111000100000001010100101000110011100011100000111011101111011001000100010010000010111110000101110101010101000010100111010100101010000110010011100110011010000001100011111001000110011010001111100101100101010011110000001110001001110000000001100001111100110000011001000110011001101000100101010110100111010000000100000010010011011101111011101011011010000111000100111000011110111011001110101001100010011101011100100101110011001010000001101010111010011100101100110101001101001011010101001111000110111101100111111000100001011111110111100110110000001110110111111000011111011010000111101110101111011110111110111000001011101010111011101111100011101000111100111111100011100111010110111000111111110111100001011110100111101001000100011010001111000011001001000101110001100000000100000010000011000011001011010010110111101110110001010000010100000101100101100101010001000010101000010100001010011100111100111010100111010111111010011001111001010111110111111111101110000111110011111111101001011111010100001111001001111110100001111101010100111100101011111011101111100101100100100110010101001101001101010111010100110100110011010100110100101101001000010010111000000110100101101000111010010000010000000101110010010111001111101001000101000010100001010000001010000100111110100000001110000010010010001001000100100001000101101001011010010110101001011010110110101101110000010101001010011101001100101010010101011010011000101000101010101000011001110110011101100110000101010010100111010011000100001010001000000110010110101010101011110010111110000110100001100100000001100010000010001100001111100111110000101110110000111110011101101110111011110000001111011010010111010101101011110011110010101101011010110100001100101111001001101110100011010110001111110100010100101001010010001101101001011011011110101010101000010111011001100010000101010101000010101000101010101000101010010001111000110011111100111101100011111000100111100010000100011010001011011010000101100010110011000010100010010100100000100001010001010100011011011011011100000101010101000100000010110010110010101101100101001110111000010110011001100001101011111110111111001010010000000100000000011011011010011010001000000010111011111000110100101101000011010010001000010011000100001000100000010000001000010001101110001101110001101111000001101001101010101010011010101100100111010010001010100101010010100000001111100111111010110001011100110111011101111010011001010110010001100011000010110010110010101110101100011001011101111010111000111100000100011101101110100101110101100011110111000101110110110110110111000010110100101110001011101100100011010110101101110000111010010010100101101010101010001111011010010000110000011100000110010110110110010010011011001110100101100010111011111001100000011001011011010100000101100101111000000000111000110110110110001110001110001110110011000000000010100010000101010010100101010001101001100110000111101100001100001100100010110001001000100001101100101101100111101100110011110011101111001111111100110100100111110011111001111000110110110100111000001100101100110100100011101011111000110110001010001100110101010110010010110111100011010001000001011101010001110110111000010100101100101100101110000110011111101000111010101001010100011010011001001111100000011110111001111101100000001011101000000011100111011101011011101100000101001010101010110010011111001011111110100011111101100100111111011001111111010011111111010000001110001001110000101110000010001101101101111100111000111011011011100001111011111100110110110110110110110111011000101111000010100011000110000111100001110111000001101001111001000111010010001101010011001100011000000110001000001101110100010111101101101111011110000101101111000001111100001000010110011100101010000101110001011101011011010000110100111001101101001100110010101100110111001100001000100101101101011110000100001110000111000010001100011111000111110001110011100011011100101111100100100111101000011100011011110100100011010000110100001101001000010101011010010101001010101101010001100100101010010101010110100001101101101001001001101000111010000110011110001100110101001010100000110110110110110010010001001000111100011100000100110000010011111010110111110100111111001010001100000011011000001110100111100000110100001010000111000011001010101011010011001001000110100100010010000010000101000001100010000101000110100001001111000100001000000010100101010011101000100100111110100001001101000110100110010111000010000011000010100010000011111110000000110000001111110111110010111011101101001100001010100001011000010000010110000101110011010101010001101011011000110001000100100001111001111011110110100111000100100000101010101000100100110101101100100011100010011100011101011110110010100001010001010010110000110011001110100101110111111100111010110010000101000001010001011001110111100011010011000111100011010001010010001101000110100011100011100110101110000001100010011110010010010000100000000000100001010000101001110101000110010111010101011111111111011001110111000111000011011001000000011010111111101111100000000001101001101101101101101100101010010100111010100001100001111011000011011001000110011011100101111001110001001110100111010100100001010101011001111100001110001001011001001100000111011000111000011001100011011001001110001000011001011110010011100100100100111110011101010001001110111101111100000011110000110011010001110100001100111000011010011001101010111010110101001111111100100110110001010100011000111011110111011101001111101011110100100100100011101101101011111111101011001100000011011100110100110110110100001110001101101001000101110101010101100001000010100010101000001000010010011100111111101001011101001100110011011100111111110011010010111000101101011011100000111011111111110000001111000011000101000101000101110001010001000011011000110110111100010001111011111011001111011000111011000100010101010100010101000100101110001110000100001010000010110000011011101111011101011011101100111000111111001001111001001000100001101101100100011100011011011100001101000011010000100110000011010011010101010100110000101011111010110101001111011010111110001011110111110001111100111011111010011111100101000110011101101000011010100001010001101000101101000111010000111010010111010111001101110111101110001101101000011101110101110111000111000001001110010011110011111110100100001010001010101011000011111001011110000100011001110110100001001011001111011101011110111100111111010000001101101111101110011101101110010001111000100010111001011010010111000101111000010011001001011100101100110011001100011111000111001010011110100101101000100101101101000011100000100100011111011010010111111000110010100101100000110111110111000011111011110100101101001011010010111010001001111100111011010010001101001111001000111001000001100111011010010110100010011110100001111100011011111110011000110100101101010110010110011001011110011011101000000101001110100010110010011001011110010101100100100011010010011010100001000000011111001111110011010100110100101101010100010111010111010111000111110011111101111100000011100010010001100001111100111111001000000100001010001110010000111000101100010100011000010111100001100100101010010111001010001100010011101010111001001001011110110111100101111010001100101101001101000011100010010111000011010011110100111101000000110011111010100110011010010101011010010101000100100001010001011000100000110000111111011000000100001010001111100001111100101111000000000101000100001011001111010011010101101011100110101100011111110000101000010101000100010101100000010001000001111001001111011100001111001111000010011110100100011100000100000011100000110110100100011110001001011101110111011101111011110000101110001001011011000001010001010100010000100001010111010111011010011101110101011011010000110100000010010101110000000111000010010001011010010110100000111111100000010000111010111001110010000010111010100101110110001101011000111111001110011101010100111000100010000010100011010001101001100100000110000010111111101100100000101101010110010000000110101111111011011111000101011001001000110000011111110110010010010111010111101011001010110010011110100111010100101001100100001110000111000011000101010101010111110001110001001110111000111011101000110101001001001110011110011001001110010011100100000101101111011011010111000001101100011101100011101101010011100111011100101111100110100110101011000101110100010011001011110010111100011100110010001100101011001000001011101010110111101110000001011101011001011010101111010010101100011101100111111111011010101011010100110000100010000100000001001110100111110011010011000101110001111100011000010000101010101100010100001010100011010001100110111001111110100010011100010011100000111011110100110110001110000001100000100100001110001001000101001100010011000110110010010011101010011000100110010000011000100010111110011100010010001011011010111000001110110100111000010111011010100010000110110100100010100010000100100010110010101010101000001100001100001110111011100101111110011101001011101000110011011000111011000011000000001100110111010000110100100011000101111011000111010101000101000001101100010010110101010100000110011010101101010100111011000110001011100100000011111011110101110111011101100111101110001111000110111011111000111110010101111101000111111011001001010000101000010011010011000101110010001100101100111110101001111101101111111011110001111110110011111110101001111110100100011111111000001111011101111110111011000111110011111001010000111000000111000011111000000000101100110001000000001110100111110100111110011110011101011111100110111100010100110110111110000101011011100011010100110111010000000110001011011011011001000111000100111011111011110101111001011011010110101101111100001011001011001011000010110011111101011100111010001111001101111000110001001010100111010010110011101010011000101110001100011111100010111110111011111101011000111010101111010111110001100011101100011001011110100100010010011001001100101100101101011011011110111110001001101100111110011010010100101010011101001000010100000100100101010110101011010011001010101101001010100010001011101111100101010001100001100001100000011111010000001000000000101010101100101100010011111001011100101100011011011011010010001001011011010010011010000110101011100110100011011011010011100000000011011001101000111001111110100010001000010100010100011110101100010011000011010001000000011111110000010010000000111111011111100010110011111001110110011000001010011100011101110100100011000010001110001001011010101011010010001011100011110101000110111100111010111100101111010011101100110010101010111000111101001100100010101010010101110110110010011100011100011100011010000001001011101001110111100010101100101000101100111011100010011010010011100011010000110110100101101100000111000110100001010001011001100000010110010110010101000110010110100111011100111011101001011010011100011011001010011101010001101100100001010000101000010001101111101101111101101111100001111110110001000001000101000001010100010100010101011110010011011110000010000101000111101101110101100101111010110111101011000001000010100010101001010001101000110100100010000101000010100000110110010101100010110101011001000000011010111111111100111010011001010010101010010101011010011001001101100110010010110010100001010001100111000100010110001001001000001000111100011110110100111111000110111100100110010101100010101011001001110110010110010110010010000011000000011111100101111011011110110111101000101000101010100100110110010110110010110110101001100111111001101110010110011101011011101011111101001000101110111011110010111110001101101011101101101101101010001101010101000110010011110011001111001011111110111100011101010011101001011101001000111100001111110101110111101011100001111101000011010110110101100011111100010010110001001011000110101101011010101001001000000001000010000010100111010010101010000110010101100100011001111001101000010010101001101001101001010010101010000001010000101000010100000010001101000101100010100100011010010001001000001111001110111001001111001010001111010011111000110111001011001001111100111110101000001010001010101010100111001101111001100111010010001101111111101111001110000010111010000001010100100100000001000011111000000110110110110001000010000110100001001011100010000001110001101101110001110101011011011001011011100111011100100110101011101000111001110000101010101010100100110111111110111011110000110010010011001010101000000110011011101000111001110001111101110011110010111111010000001111011110111110111000111100010100110110010110000101100001000011001101010101010000111000100111000010110111111001101111001101111101101111100010110100101110111100000000110000111101101111010100001110100011110011001110001110011001111110011011100011100010110010111100000000011000010100010101001110111101111100001011110110111000111111010111011011001000111101101101001000000100101111111000111001001011100110010010100010001101011100110111010001100101011001000110001010011110100011111101101111111011011001110100011110101101100011000110010011101000011111001010001001111100110110101000001110001100101110111000010111010110100101101101010100101010110101001010100001100111011001101110001010010100101010010101010100011100010010111000010000001000001011111100010110011000010110000100101101101101100010100000101100010010001011011110111011000101000101100101010001101101101101100100101000110011101001110001001110100110110011000010011101001101100111000101010110101000110010001111100110000111110001000000100000110000000001101101101101101000101010110100111010101001010101101010110100100111010100100101110101000010010100000101010100001011000000100100000110111010111010111101100000011110110100110101010000111100101111110010100100101001011100000100001000010101011101100110010111000111000111000001110001000011101011111010111101001001010000100000010000001110101001000110100001000000100100011010011011011011011101111000110110001010001110000010110010101010111101011101110000101010000100100011100000001101101100100010101010101011111100010111010110010101000110010110010111000001111110101111000000001100000110111111101111000011101101111110110111111011010100111100000111101111011111000001000111110010110010110011110010101111011111101011000101101001001011101111011000111100010001011000011100011011010100100000001010001010101111100010100111010011101010000100000110000011011001010110001011010101100100000001101011111110110001000000100101001110101000010011100110010111001100100101000100101010010101101010100100100111010100110100110111100011100000010001000001011101110111010101111010001010001010001010100100100010010001011010011110101100111110001111101011011100100100110101011111011000010100011011010000011000000101111111011111100111010011111010100111010000001101101111101110001101110110010110111101110001011011100110101011101010111010010001010000100111010011000001011101010101000001010011101010110101000010001101000000100000000111000011111000011111000011001000000100000110000001011000000010000101001110111011000010100011010001010111101001101100000111010011111110101001101101101101110000101010001100101100100100011010010001011010000111101100001111011000111110101111001110011111110100011110100110011110010111111110000111110100010010011011001100100110000111110110111111101110011111100000001111001100111100111011100010100000001011000011100011010011011001000001100001010000010001010001010000000101110100001110110111011011101001010101010101110111000100011101000101010101010100000010101011010010000001101101010001000000110110110110101010001101101010001110111110101101011011100010110110101101010011011101111011110011011110100111001011111001011111101000000111010010111010110110010100010101001010101011001001000100100000101100000101001110100010110100010100101010100010010011111101001111111111000001111011111100111010101110001111101000000011000010101101001100110000001011110110111001001101010111010010110011110011001110110010111100101000110000101100001111011101000101111001011111011000001000110000111110010110001101010011010100110100110010111110110110110110110100001011101010111100110000010010010101001001110100010011000101111011000111010010001110100101110110001100011100111100111111100100111100101000111001011111001011111010011001100111011001110110100100001101101000010010011001011110010111100100000011000011111001111110001111100101010101100011010010110100011100110100100000010000001000100000001000010000001110001101001101100011111001100001100000011111101111110111111001000010100001010000100001111101000000011111001110100000111001010011001001110001001110100101011010100001010001101000011010101000110100110100110100001111100110001000101000101100101010101100001010001010101011000100001110000011000011000001000010010001000011110000000000010011010011010101010100011011011010101010000010101010110010110011101011100100110100001111001010011100111101110101110010000010000101000111101010010101101111010110101001011110111010111001110001010100001001000101000100101001011110101100001101000011011000110110100101110101011100001101001011101010001111101010111011100111000100001110110011011100110011011000111000100001010000010110010111010111000100001101100001010100011001011011000110100110011010100001000001011111110000000011000011110000011101100110011011110011011110011011110100110000101100001011000001000101110110000101000010000111000011100000000101001110101001010100001000111100011001010010101100010101100011000010100101011000000110101010110000110001010001001010110000111001000000100000000101010010100101010010101001010110011101001100110100010110010000000110101111010110101010010000111001101100101010010101001010100011101010111001001010110100111100111100100101110010011101001000100110010010111001100001010101101010101101000011010011001101010100101010110100111010011001000100100010110001100010010011101010011010010001000000100000110000100010000001000000100000100011111101111110111111111111101011011001101110011001001010010100100011011011100011011001000010100010010001100010110110101101101011100000110001011100010111101011100100100010010001001000001101010011010100110100100001011001010101011100100011010001001000110001000100100001010001100001011101111100111110000101010101100101100111010111100100010111011011011100001001111101000110100000011100010111100100011100011100101101011001000100100000110110101110110100110110100000111110011111001111100010101001010101101001100100100110010101001011001101000111010011100101000110100101101010010011000010100101010010101000000101001010100011001111001000110100011110110100001011100010111001101110010011001010110011111100111000101000110100001010010000111110011111110000100010000001000000011000001010101011100101001000010010001110100111010010110101110001011011010001000001100001111100101010001001010100010110000101000101010100100011100011100011011000101000101010100000011100011100010110110101110001000101000110000010100001110000111110000101101111110010011111001011111101111000011110010101111101101011111010110001011111111000000110110001001110111000111011010111011100000110110111110110111110000000010000011000010100011000110100101101000011001101001110101111110101001110011110010111000101101111011010100011100011010011100001001000100100010110100001101100001101100011101100100011101101011110111001111100000001111001000101100100101101100110011111101010011111100000001001101101000110011100011001111111010001111001101001111101100111111010111111110101010011000100111010111111011000001100011011001010110011110010100001010001101001000101101011011100010111110001001101100110010011000001010001000011001000111110010111011111100101000010100001001111001001111010010111000001011101100010000010000010100010111000101110111110010111000111110010100010101001010010101000110100010001111110110001000000000101000001010000100100111010001110100110111011001100000001001010001010000101000010011111001100000100000010100000111110011111010000011010111110001001101110001010101010101011000010100010100010100101011110110001011100001001101011001001101100000001110001110000010100011100011011000100101111001111101011110101011000001111011100010001101011010111111001100001111010100110011111011100011110111001110000000100100011011000101000001110001110100100000001111010000100000011011011100011100000100001001010010001101001110000000101010101100101010111010111001001001000011100011101111101111010100110010110101010100000101000101100100000100000010000100111111001011111010001111011110100110110011110110100110111000001101100111100001111000001001100001011000001101110100011101110001110111000111011101100110100011101001010011010011110100101110001101110001100010001101011010010110101001110011001110100011110100100011100010011100001110000000010110100100011001110101101001000111000100010101100101011000011111010111101001001000011101011011001000001000001010110001001001111110001001010010010100101010010101001000100000010110010100111011100001011001000000011010101011000000100101010100011010010101000100100110110011001001010001101001011010010110011110010010101001001110101000010011111001110100110100011001011001011010001010011101000101110111010010100011001010101010110010100000101100101010111110001011010010111010101110010010101000110011010010001001111101001010100100011001011110010111100101000000001010000110110001110110010110110100111111101011010011100101101010101101101100001010001110111001101110001011100100110001001100010011101011000100101010010011001011001110101011110100111110101000001011001010101010000101111101011110010111011000101010101100101100001010101011001010100010010111101110100011100010010101001010100101000110010111100111111010001001100100011001011110011000011001010110010001100101100111100000011101110101011101100100110110011111001111001101001111010101110101010011000111110011101100110000110011111101000110011000010101001001110011001001010101011010011011000100101110001000000110110100101001001100101011010001110011010001101101101101101100011000011111110001000001101101100101101100010101010101011000000101010101010111110000101000101000110010001001010010000011011011011000001100010000011000000011101111010000011100101010111011001101001100001001011100010110011110011010101110001111010110111011001010111010000111100010000100001101010001010001000001111011011011110110101111100011100101111111011110110111100001011110010111001100011100110100101100100111100011100110101001100110111000101000110010110110101000010000111000011100011000111100011111110001011111011010100010100010101100000000011000100000101100000100000110000000110000011101001111101000111100110100011111001111110111111001101000111010011110100010011110011111111001011111110110000011100010111100101111101001000110100001001010111110101110001101010101010110100010011101010001101001000010100010110010110000101100101100111110001010100101010110100000011010100110100111101001000100110010010101001011000001001011010001000100100010010001010001100001111101000001000100100010010001100001100010000110001111111000010100010000010000101000111011010011011101010100111010100011001001001010100110010010110001101010101001010011001010101101001110100110010000011000010011101011010100111010001011001010101011101111011000111110111000101001010111001001111010110000010100011110010010100100000010100011110111011000101000011010101011101101110011011000100001010001011000010100010100011101001110010000010100101001011101101110101001110011101101101100011000011101010100000111111011100010010111011010010101100101010001010001010110110000011110011111101001110101100000011000010101000101000101010000010000101010001101101110001100100011100000110110001010101110001110101001101110000000010010111011111111011110101110011011100110111011001101101001101101011101101110011101110011110110111111011010000111000011111000010111000011001101000110010011001100001110101011110101001110100100011100011011100101111101001000100000010001101000100001110110101111000000111011010100110111111101000011011101100111010011110001001110101010010000011000100100001000111001100111001100111010001001110111001111000100111011010000100000001100010000001101011111100011110001010001110110011010110101101110101011000111110011010010110000110110110011010100101100100000101101011111100111100110000000110100111000111000110110010100011010001101000100100101010011001101010100110101001101001011010000001001011100100111010100001001101100111010011100001101101101001101110101111011101010000100110110110110111000000010010101100001011101111100111111000111000100110101010000010000000110000111101100111101101000010011001001110100101000110010001100011111101100000100010010001001000101001101001111010011110100100010110110101110001011101011111100011011100111101011110010100011110010100110011011101000010100001010000000100001010001000001101100101101101001101101000001001011011011011001010101011001101001100110001001110101011110101000010000111000010100000100100011110110100100100000010111010000101101010111000101011000110100111101010110011000011100010111100101111101010000010100011010011100001111011011011110001011111011010100101111101101101101011101000111110100101111101000011111010111001100010111000110110011010010100111010101011011000111000001000000101010001010110101111110100010111001110001111011100110000111010110010111011000001011010010110110101111010001011101111100110000001010101010101010100010111010111011111101110100111101111100010100010000001010101010001011000101001010101000111000001011001010101010100011000011111001011100010010100001010000011011011011011100000101000111101001100110101001000101011101000100000100101110101001011000100010101101111110111101110110101111011011111100000100111001000111000101111101000100010010110100101000001000010010111000010111011101111001100000100101001010101011010100001011110111011000011000010001011011010111001101111100010011101001100100101100111010100111010001111001011001100110111001111110011010011111110100111111001101111110010010011100110011100111011100111100110100001100100111010000001001110101000001100100110011101100111111001110001001000100011110001110010011011010000101000000101000010100011001111001000011100001101110110100101101100100111110011111001111000111110011000010111000111111011111110001100010001011000010100001100100000110001001000110001001010100101011010100001010010101001010100100000010100010100001001011110100111101001000000100000000101110111111100000000010000001000000101110111110011111100010111011000011111101110101000111100010100000111011100111001011110000000010101010001010110001011101010111011000010110011100100001111010011010110100011100011011000001101001101101101100011011011011010010001000000101000001010001111000111111101010000111101100110101111110101011000111011101010011100010010110110111100100110000001000110110001011001111001010011010111101110101010011110011101110000000110110110110001010101010001110100000010110101110010101010110100001101101101001110101011100100101010111010101101101011100000110111000110110101110111010001101111101101111111101111100001111100110001000001001000010011111101100000010110011111001001001000111101101001000101001000101100011010001100011001011110010111100110000110110000110110000011000001101000011001101100101000110001101001000110001010011011010011011010011000011001001010100110110010110011010101100100110010010001010101100001011000111001011111001111111010000001110111000111011010011101101001010111110001101111001010100111010010101010000000001001001000000100000101110110011011010111011011011011011011000101011010111101001011101010111011110001110101011010011001101010000101010110101011010101101100101010110000111111111100111101000000000110100110110110110110110010100001010000100111100100110010011011001010001101010111010100110100000010010011101010011010100001001100100110010011010001101001100101100110101111100000000000011001011000110100111010000010010100100110110100110110101110110100001011011110111010101110110011100011011100010111110011010011010100100101011001110001111010011111000101101010000111000100111011101011101111010001010011001001110001110011010101110100111101000100010100010101010110001100111011001100110010100010001001000100110111001011110111011100101111010001111010100000000001101001110100000011100001011100011010011001011001001010011101001010100100010001011000100100011000101111011011111010111111001011010110110111101101000010010101101010111010101001101000111010100110101000011100111011101001111101010100101111001011101010111011001101101101101101001101100110010001001000100100001100110111011110111100110111010001111101111011111100000111100110000101110101011010010110111001011110111011000110110110001111100011111111001011111110011100011000110110001001101000000010010100001010110101111110100011011001101101000011101111010000100010101010101000100001110100100101000011010000100101111000101011010100011100011101011001000001111001000000111101111111011101010101000101000101100101010001000010100010110001001011100101010010010010011001001100110101010010111001101110001011110001110110011000011010011110110001110100010001000010100010000111010111001000000101010100011101010101100100111010101010101010110000101010111101111101011101101011011011010110110001100001011011001011011011000010101010001101100100011011000011000001101111100000000111000011110100101111001101111110111100011001111110011101100101100110011001101001111010011001111101100111111011000111110111000011100100111100100011100101000110011001100110111001111000100001011101111100111010101100111110101010010101001100010111011000011111100010110010111010110001101001111010101110101001010111110100001101010001010101101010110101010001111111000000100000100010111011111001000001010011101001010011100010110100101101001000111000101000100101000001010000100111010010100000000111000001100101100110101010001100101100101100100011100010000100110101111101100001100110001010001010001010101111010011010111000010011101011001101110110011001011000001011100100101011010110011010000010110000000001010001000101011101001010110000001000010000101000010101011010101011010011101000000011010011110111000110110010101101101010000010011000010010001111011111111011111001110111111010110110110110110111101100010100101100011011011011000101100101010101010001010100010101011110011100011101010101110000011001101010110101010010000010110001000001001011011010110100101111100011000010110110001110000110011000011110110010110110001001011101110111010100100000111011010111100001111100000100110000111100001111011010000111000110111001000111001111001001100100100111010010000100101110001010100111010000111010010111010001001110110100110111111110111110001110110101111000000110111101001111001100111100111011110011010010001111011010010111011001110101101100010011000111001000010100000110000000011100001111100000111011110000111000101111000111111001111001000001100000101011000100010010001001000010001100111011010000110100100010100111010100101001100011111001011101111100010001001000011100010000100100110010011001010000111110011000010100000110000111110011111100010010110100110010001010101100001111110010110111101101001001000000100001010001110110011001001110010111011111001100000101010110101011010100011101001110100101101011001011010010010110011111100110110010000000110100110110110110110110010100101010010101000000100100110010101101010100110100111101000111001111001001010100101011010101001001110100111010011100001110001101001101001111010111010101110010110001001000001110010111100110100010001110101011011011010101110100010100010000011010000110011111100110000101110111011110110111110001011011110111001101110100011111100001111111000001111001100000110000101100111111000111111100000101111110010101010110011010101000110011010101101010100011000011000100000000110100111101001011010001001100001011011000111011001000100000010000001000000111101010101010101110010011011100011100011100001010011101001110100110001110000010010011001001110001111100100000100100010110101100011100110010001100101111001000001011011010110100101101100011011011111011100111011100100111100110111110100111111010010001100010111001010110011110011010010110101011001100001000100100011110010000011101011111001111110011110011100110011100110111101000000110011111101001011010101001100111111001110110100110011001000111111110111111010010001001111101000101101100000001110111011001000010011010011011000001101100001000110100001000010011101011001110110010100000001111011000101001111000100101101100010110011111010000000111101010011110110001101110101111001101011001001010101011001000001001011100101111010010001110100101110100001110011100010001111110111001101101010001100010000000101100001010001011001011101110110011011111010010101010101011101001110010101001101011100000010111010100110101111011101111110101101101001101101001101100110011101000011101000111100110100111010010111010100111001101001100010011101001011101000100111000111111001011111001111001100111111010001100101000101000110101010111000010011101001111101001100010101011111110000000010101000110110100000101010010100011001111000100101000101000000100110010010101001100000111111100000001100000100000001011101011100010100010101010100000101110101000100000100000010000101000101001000001100010010000110001111110111111011111100010100010010101010011001001110010011010000001101010011010100110101000010101011010011101000100101001010011111001011001000000100010010001110001010001010101111110001000010100010101001000000100000101110100111011100010011100011100011101110000111000001101110111100011001000100001111001110101101100000101101011000000110100100111010100001010110110011110101111001000101100001100010011010010010000101000101000001110001101000101011111001101010111101010110111100011000100000010100011110101001000000010111000001001011011011100000101110100001111100001010101011001010100011010011110110101001110011110110100111101100001001110011010101010000101100000010100010101001000101100011010001100011011001011000011110000110011100000111011100011011101000;

reg clk=1'b1;
always #10 clk = ~clk;

reg         ivalid = 1'b0;
wire        iready;
reg         ibit= 1'b0;
wire        ovalid;
wire  [7:0] obyte;
wire        raw_format;
wire        end_stream;

task automatic test_codelen_tree_build(input logic [BITSTREAMLEN-1:0] bitstream);
    @(posedge clk) #1
    ivalid <= 1'b0;
    ibit<= 1'b0;
    for(int ii=BITSTREAMLEN-1; ii>=0;) begin
        @(posedge clk) #1
        ivalid <= 1'b1;
        ibit<= bitstream[ii];
        if(iready) ii--;
        //@(posedge clk) #1
        //ivalid <= 1'b0;
        //ibit<= 1'b0;
    end
    @(posedge clk) #1
    ivalid <= 1'b0;
    ibit<= 1'b0;
endtask

initial begin
    test_codelen_tree_build(bitstream);
end

always @ (posedge clk)
    if(ovalid)
        $write("%1d ", obyte);

huffman_inflate dut(
    .rst        ( 1'b0       ),
    .clk        ( clk        ),
    .ivalid     ( ivalid     ),
    .iready     ( iready     ),
    .ibit       ( ibit       ),
    .ovalid     ( ovalid     ),
    .obyte      ( obyte      ),
    .raw_format ( raw_format ),
    .end_stream ( end_stream )
);

endmodule




























module tb_huffman_decode_symbol();

localparam BITSTREAMLEN = 327;

localparam NUMCODES = 19;
localparam CODEBITS = 3;
localparam BITLENGTH= 7;
localparam OUTWIDTH = 6;

function automatic integer clogb2(input integer val);
    for(clogb2=0; val>0; clogb2=clogb2+1) val = val>>1;
endfunction

reg clk=1'b1;
always #10 clk = ~clk;

reg                   ien = 1'b0;
reg                   ibit= 1'b0;
wire                  oen;
wire [OUTWIDTH-1:0]   ocode;

reg         wren = 1'b0;
reg  [31:0] wraddr = 0;
reg  [31:0] wrdata = 0;
reg         run = 1'b0;
wire        done;

wire [clogb2(2*NUMCODES-1)-1:0] rdaddr;
wire [            OUTWIDTH-1:0] rddata;

wire [31:0] data1 [NUMCODES] = {3,5,6,5,0,4,5,4,3,3,4,3,4,5,5,0,6,5,5};

logic [BITSTREAMLEN-1:0] bitstream = 'b111110110011000100011010001010010101010100111101110101010101101110110001011000000110110000111110101111111111101100011101011111101111010111111011100011000000110110000000110110110000111010101000100110011000100010001100111100001001111011000100100110101001010000110100101010100101010010010100010010100010010011001010110011100011000;

huffman_decode_symbol #(
    .NUMCODES( NUMCODES ),
    .CODEBITS( CODEBITS ),
    .BITLENGTH(BITLENGTH),
    .OUTWIDTH( OUTWIDTH )
) dut2 (
    .rst     ( 1'b0     ),
    .clk     ( clk      ),
    .ien     ( ien      ),
    .ibit    ( ibit     ),
    .oen     ( oen      ),
    .ocode   ( ocode    ),
    .rdaddr  ( rdaddr   ),
    .rddata  ( rddata   )
);

huffman_build #(
    .NUMCODES( NUMCODES ),
    .CODEBITS( CODEBITS ),
    .BITLENGTH(BITLENGTH),
    .OUTWIDTH( OUTWIDTH )
) dut1 (
    .clk     ( clk      ),
    .wren    ( wren     ),
    .wraddr  ( wraddr   ),
    .wrdata  ( wrdata   ),
    .run     ( run      ),
    .done    ( done     ),
    .rdaddr  ( rdaddr   ),
    .rddata  ( rddata   )
);

task automatic test_huffman_decode_symbol(input logic [BITSTREAMLEN-1:0] bitstream);
    @(posedge clk) #1
    ien <= 1'b0;
    ibit<= 1'b0;
    for(int ii=BITSTREAMLEN-1; ii>=0; ii--) begin
        @(posedge clk) #1
        ien <= 1'b1;
        ibit<= bitstream[ii];
        @(posedge clk) #1
        ien <= 1'b0;
        ibit<= 1'b0;
    end
    @(posedge clk) #1
    ien <= 1'b0;
    ibit<= 1'b0;
endtask

task automatic test_huffman_build(input logic [31:0] data [NUMCODES]);
    @(posedge clk) #1
    run <= 1'b0;
    wren<= 1'b0;
    for(int ii=0; ii<NUMCODES; ii++) begin
        @(posedge clk) #1
        wren = 1'b1; wraddr = ii; wrdata = data[ii];
    end
    @(posedge clk) #1
    wren = 1'b0; wraddr = 0; wrdata = 0;
    @(posedge clk) #1
    run  = 1'b1;
    @(posedge done)
    @(posedge clk) #1
    @(posedge clk) #1
    run  = 1'b0;
endtask

initial begin
    test_huffman_build(data1);
    test_huffman_decode_symbol(bitstream);
end

always @ (posedge clk)
    if(oen)
        $write("%d ", ocode);

endmodule























module tb_huffman_build();

localparam NUMCODES = 19;
localparam CODEBITS = 3;
localparam BITLENGTH= 7;
localparam OUTWIDTH = 10;

reg clk=1'b1;
always #10 clk = ~clk;

reg         wren = 1'b0;
reg  [31:0] wraddr = 0;
reg  [31:0] wrdata = 0;
reg         run = 1'b0;
wire        done;
reg  [31:0] rdaddr = 0;
wire [OUTWIDTH-1:0] rddata;

wire [31:0] data1 [NUMCODES] = {3,5,6,5,0,4,5,4,3,3,4,3,4,5,5,0,6,5,5};
wire [31:0] data2 [NUMCODES] = {3,6,0,7,7,5,7,5,4,4,4,3,3,2,0,0,7,4,6};
wire [31:0] data3 [NUMCODES] = {3,6,7,6,6,5,6,5,5,4,3,3,4,2,7,0,0,4,6};
wire [31:0] data4 [NUMCODES] = {2,7,0,7,7,6,7,5,5,4,5,3,3,2,7,0,0,5,7};
wire [31:0] data5 [NUMCODES] = {2,6,0,0,7,6,7,6,6,5,5,3,2,3,5,0,7,4,7};
wire [31:0] data6 [NUMCODES] = {2,6,0,0,7,6,6,6,6,6,4,4,3,2,4,0,6,4,7};
wire [31:0] data7 [NUMCODES] = {3,6,0,0,6,7,5,6,5,4,4,3,3,2,4,0,0,4,7};
wire [31:0] data8 [NUMCODES] = {2,6,0,0,6,6,6,5,5,4,4,4,3,2,7,0,6,5,7};

huffman_build #(
    .NUMCODES( NUMCODES ),
    .CODEBITS( CODEBITS ),
    .BITLENGTH(BITLENGTH),
    .OUTWIDTH( OUTWIDTH )
) dut (
    .clk     ( clk      ),
    .wren    ( wren     ),
    .wraddr  ( wraddr   ),
    .wrdata  ( wrdata   ),
    .run     ( run      ),
    .done    ( done     ),
    .rdaddr  ( rdaddr   ),
    .rddata  ( rddata   )
);

task automatic test_huffman_build(input logic [31:0] data [NUMCODES]);
    @(posedge clk) #1
    run <= 1'b0;
    wren<= 1'b0;
    for(int ii=0; ii<NUMCODES; ii++) begin
        @(posedge clk) #1
        wren = 1'b1; wraddr = ii; wrdata = data[ii];
    end
    @(posedge clk) #1
    wren = 1'b0; wraddr = 0; wrdata = 0;
    @(posedge clk) #1
    run  = 1'b1;
    @(posedge done)
    for(int ii=0; ii<NUMCODES*2; ii++) begin
        @(posedge clk) #1
        rdaddr = ii;
        @(posedge clk) #1
        $write("%d,", rddata);
    end
    $write("\n");
    @(posedge clk) #1
    run  = 1'b0;
endtask

initial begin
    test_huffman_build(data1);
    test_huffman_build(data2);
    test_huffman_build(data3);
    test_huffman_build(data4);
    test_huffman_build(data5);
    test_huffman_build(data6);
    test_huffman_build(data7);
    test_huffman_build(data8);
end

endmodule
